"Normal string"
"Weird "" string"
"even weirder " "string"
