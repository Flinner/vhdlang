-- This is a comment





-- This is another comment
